module controller(rst, clk, imHeight, imWidth, imAddr)

input logic rst, clk;
input logic [7:0] imHeight, imWidth;
output logic imAddr;

endmodule